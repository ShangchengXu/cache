interface list_ctrl_interface_inner;




endinterface