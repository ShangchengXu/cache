class memory;
static   bit [31:0] mem [4096];
endclass