interface rd_ctrl_interface_inner;




endinterface