interface cache_ctrl_interface_inner;




endinterface