interface wr_ctrl_interface_inner;




endinterface