interface ro_cache_ctrl_interface_inner;




endinterface