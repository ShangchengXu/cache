class memory;
static   bit [31:0] mem [4096];
static   bit [31:0] mem_model [4096];
endclass