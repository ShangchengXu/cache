interface mem_ctrl_interface_inner;




endinterface